library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity D_TRIGGER_ACCESS is
    Port ( D, CLOCK, CE : in  STD_LOGIC;
           Q, nQ : out  STD_LOGIC);
end D_TRIGGER_ACCESS;

architecture Behavioral of D_TRIGGER_ACCESS is
	signal out_value: std_logic;
begin
	p1: process(CLOCK, CE)
	begin
		if CE = '1' then
			if (CLOCK'EVENT and CLOCK = '1') then
				out_value <= D;
			end if;
		end if;
		
	end process;

	Q <= out_value;
	nQ <= not out_value;

end Behavioral;

