library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity RS_TRIGGER is
    Port ( R, S, CLOCK : in  STD_LOGIC;
           Q, nQ : out  STD_LOGIC);
end RS_TRIGGER;

architecture Behavioral of RS_TRIGGER is
	signal out_value: std_logic;
begin
	p1: process(CLOCK)
	begin
		if (CLOCK'EVENT and CLOCK = '1') then
			if (R = '0' and S = '1') then
				out_value <= '0';
			elsif (R = '1' and S = '0') then
				out_value <= '1';
			elsif (R = '1' and S = '1') then
				out_value <= 'Z';
			end if;
		end if;
	end process;

	Q <= out_value;
	nQ <= not out_value;

end Behavioral;
